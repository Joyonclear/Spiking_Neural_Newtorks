`ifndef PARAMETER_NEURON_VH
`define PARAMETER_NEURON_VH

`define DATA_LENGTH 32
`define MAX_THRESHOLD_VOLTAGE	4080218931	//2**32*0.95
`define MIN_THRESHOLD_VOLTAGE	3650722201	//2**32*0.85
`define MAX_RESTING_VOLTAGE		 644245094	//2**32*0.15
`define MIN_RESTING_VOLTAGE		 214748364	//2**32*0.05

`define RESTING_CONTRIBUTION	   8589935	//2**32*0.1*0.02
`define THRESHOLD_CONTRIBUTION	   8589935	//2**32*0.1*0.02

`define RESTING_DECAY				 42950	//2**32*0.1*0.0001
`define THRESHOLD_GROWTH			 42950	//2**32*0.1*0.0001

`define TAU						1024

`endif
