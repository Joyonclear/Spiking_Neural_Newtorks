//############################################################################
//## Neuron design Num.02 => LLIF model
//## Target device : Xilinx XCZU9EG-FFVB1156AAZ-1e
//## 
//## designed by Huiseong Noh
//## File created : 2021-03-13
//## Last edit : 2021-03-13
//############################################################################

//############################################################################
//## Info.
//## test bench for 02 LIF model
//############################################################################

`timescale 1ns / 1ps

module test_bench;
		reg clk;
		reg[31:0] in;
		reg rst;

always
	#5 clk = ~clk;

initial begin
	clk = 0;
	in	= 0;
	rst = 1;

# 5000
# 10
	rst = 0;
	in = 900000000;
# 10
	in = 0;
# 60001
	in = 900000000;
# 10
	in = 0;
# 50002
	in = 990000000;
# 10
	in = 0;
# 45001
	in = 900000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;
# 35001
	in = 1000000000;
# 10
	in = 0;

# 30000
	in = 1100000000;
# 10
	in = 0;
# 30004
	in = 1200000000;
# 10
	in = 0;
# 25003
	in = 1300000000;
# 10
	in = 0;
# 25001
	in = 1400000000;
# 10
	in = 0;
# 25000
	in = 1590000000;
# 10
	in = 0;
# 20000
	in = 800000000;
# 10
	in = 0;
# 20000
	in = 800000000;
# 10
	in = 0;
# 20000
	in = 800000000;
# 10
	in = 0;
# 5000
$finish;
end


neuron02_LIF u0(
		.i_clk(clk),
		.i_rst(rst),
		.i_spike(in),
        .o_spike_lid(),
		.o_spike_exd()
	 );
    
endmodule
